module gates(input in, output out);
    assign out = ~in;
endmodule
